`define DWIDTH 8
`define FIFO_DEPTH 16
`define PTR_WIDTH 5
`define MARGIN 31
`define PERIOD  10.0
`define NUM_STRESS_LOOPS 100
`define NUM_OPERATIONS 50
